`timescale 1ps/1ps  

module exp_interface (clock, reset_n, );
    
endmodule: interface